package pack;
  
 import uvm_pkg::*;
`include "uvm_macros.svh"
`include "Transaction.svh"
`include "Sequencer.svh"
`include "Driver.svh"
`include "Monitor.svh"
`include "agent_config.svh"
`include "Agent.svh"
`include "Scoreboard.svh"
`include "env_config.svh"
`include "Environment.svh"
`include "randSeq.svh"
`include "Sequence.svh"
`include "personIn.svh"
`include "personOut.svh"
`include "test.svh"
 
endpackage:pack
   