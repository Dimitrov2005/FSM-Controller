interface iface (input logic clk, rst);
   bit x1, x2;
   bit cs;
endinterface // iface
